module uc(output wire s_inc, s_inm, we, wez, output wire[2:0] AluOp, input wire, clk, zero, input wire[5:0] Opcode);

endmodule